module SR_NAND_test ;
    wire Q , Qn ;
    reg R , S , clk ;

    SR_NAND aa(.q(Q),.qn(Qn),.r(R),.s(S),.clk(clk));
    initial begin
    #0 clk = 1 ; S = 0 ; R = 1 ; 
    #5 clk = 0 ; S = 0 ; R = 1 ; 
    #5 clk = 1 ; S = 1 ; R = 0 ; 
    #5 clk = 0 ; S = 1 ; R = 0 ; 
    #5 clk = 1 ; S = 1 ; R = 1 ; 
    #5 clk = 0 ; S = 1 ; R = 0 ; 
    #5 clk = 1 ; S = 0 ; R = 0 ; 
    end
    
    initial begin
    $display("HEM -- 202053007 -- SR Latch NAND-- Structural");
    $monitor ( "\nClock = %b, S = %b, R = %b, Q = %b, Q' = %b, time = %2d",clk,S,R,Q,Qn,$time) ;
    end
endmodule

module SR_NAND (q,qn,r,s,clk);
    output q,qn;
    input r,s,clk;
    wire r1,s1;
    nand na1(s1,s,clk);
    nand na2(r1,r,clk);
    nand n1 (q,s,qn);
    nand n2 (qn,r,q);
endmodule
